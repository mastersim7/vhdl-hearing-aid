-- Description:
-- filterblock_main.vhd
-- Author: Shwan Ciyako,Anandhavel Sakthivel
-- It is still in the implementation phase. 
-- This files adds needed components together to make a filterbank, you are welcome to make changes but make shure to update the whole chain of files that will be affected

-- 2011-03-30, Mathias Lundell
-- Works essentially in the same way. There is still a simulation error which
-- I believe is constrained to simulation and not implementation on fpga.
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_signed.ALL;
USE work.EQ_data_type.ALL;

ENTITY filterblock_main IS
	  GENERIC(
            NUM_BITS_OUT : NATURAL ;
            NUM_OF_SAMPLES : NATURAL ;
            NUM_OF_COEFFS : NATURAL ;
            NUM_OF_BANDS: NATURAL );
    PORT( 
            clk     : IN STD_LOGIC;
            sample1 : IN sample;            
            sample2 : IN sample;
            updated : IN STD_LOGIC; 
            Q       : OUT Multi_Result_array;
            done    : OUT STD_LOGIC;
            next_sample : OUT STD_LOGIC;
            sample_nr : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END filterblock_main;

ARCHITECTURE  filterblock_main_arch OF filterblock_main IS 
-- constants 
CONSTANT CO:taps_type:=
(("0000000101110","0000000110010","0000000110101","0000000111001","0000000111100","0000001000000","0000001000011","0000001000111","0000001001010","0000001001101","0000001010000","0000001010011","0000001010110","0000001011001","0000001011011","0000001011101","0000001011111","0000001100001","0000001100011","0000001100100","0000001100101","0000001100110","0000001100111","0000001101000","0000001101000","0000001101000","0000001101000","0000001100111","0000001100110","0000001100101","0000001100100","0000001100011","0000001100001","0000001011111","0000001011101","0000001011011","0000001011001","0000001010110","0000001010011","0000001010000","0000001001101","0000001001010","0000001000111","0000001000011","0000001000000","0000000111100","0000000111001","0000000110101","0000000110010","0000000101110"),
("0000000100101","0000000101001","0000000101110","0000000110011","0000000111000","0000000111101","0000001000010","0000001000111","0000001001100","0000001010001","0000001010110","0000001011011","0000001100000","0000001100100","0000001101000","0000001101100","0000001110000","0000001110011","0000001110110","0000001111001","0000001111011","0000001111101","0000001111110","0000001111111","0000010000000","0000010000000","0000001111111","0000001111110","0000001111101","0000001111011","0000001111001","0000001110110","0000001110011","0000001110000","0000001101100","0000001101000","0000001100100","0000001100000","0000001011011","0000001010110","0000001010001","0000001001100","0000001000111","0000001000010","0000000111101","0000000111000","0000000110011","0000000101110","0000000101001","0000000100101"),
("1111111101011","1111111110000","1111111110111","1111111111111","0000000000111","0000000010001","0000000011011","0000000100111","0000000110011","0000000111111","0000001001100","0000001011001","0000001100111","0000001110100","0000010000000","0000010001101","0000010011000","0000010100011","0000010101101","0000010110110","0000010111101","0000011000011","0000011001000","0000011001011","0000011001101","0000011001101","0000011001011","0000011001000","0000011000011","0000010111101","0000010110110","0000010101101","0000010100011","0000010011000","0000010001101","0000010000000","0000001110100","0000001100111","0000001011001","0000001001100","0000000111111","0000000110011","0000000100111","0000000011011","0000000010001","0000000000111","1111111111111","1111111110111","1111111110000","1111111101011"),
("1111110111100","1111110110000","1111110100110","1111110011101","1111110010110","1111110010010","1111110010000","1111110010010","1111110011000","1111110100010","1111110101111","1111111000000","1111111010100","1111111101011","0000000000100","0000000011111","0000000111011","0000001010111","0000001110001","0000010001010","0000010100000","0000010110011","0000011000010","0000011001100","0000011010001","0000011010001","0000011001100","0000011000010","0000010110011","0000010100000","0000010001010","0000001110001","0000001010111","0000000111011","0000000011111","0000000000100","1111111101011","1111111010100","1111111000000","1111110101111","1111110100010","1111110011000","1111110010010","1111110010000","1111110010010","1111110010110","1111110011101","1111110100110","1111110110000","1111110111100"),
("0000000010101","0000000100010","0000000110000","0000000111101","0000001000101","0000001000111","0000000111111","0000000101101","0000000010001","1111111101101","1111111000010","1111110010111","1111101101111","1111101010000","1111100111111","1111100111111","1111101010011","1111101111010","1111110110001","1111111110100","0000000111100","0000010000011","0000010111111","0000011101100","0000100000100","0000100000100","0000011101100","0000010111111","0000010000011","0000000111100","1111111110100","1111110110001","1111101111010","1111101010011","1111100111111","1111100111111","1111101010000","1111101101111","1111110010111","1111111000010","1111111101101","0000000010001","0000000101101","0000000111111","0000001000111","0000001000101","0000000111101","0000000110000","0000000100010","0000000010101"),
("0000000001110","1111111110000","1111111010011","1111111000101","1111111001101","1111111100111","0000000000100","0000000010011","0000000001011","1111111110100","1111111100111","1111111111001","0000000110011","0000010000010","0000010111011","0000010110010","0000001001111","1111110100100","1111011101101","1111001111001","1111010001001","1111100101011","0000000101110","0000100110110","0000111011011","0000111011011","0000100110110","0000000101110","1111100101011","1111010001001","1111001111001","1111011101101","1111110100100","0000001001111","0000010110010","0000010111011","0000010000010","0000000110011","1111111111001","1111111100111","1111111110100","0000000001011","0000000010011","0000000000100","1111111100111","1111111001101","1111111000101","1111111010011","1111111110000","0000000001110"),
("0000000001000","1111111110111","0000000000111","0000000110111","0000000101001","1111111010011","1111110110101","1111111110101","0000000010010","1111111101100","0000000001111","0000001111101","0000001011101","1111110011000","1111101010010","1111111100110","0000000101101","1111111001100","0000000101000","0000101101100","0000100101101","1111001111010","1110011001010","1111101001001","0001100110111","0001100110111","1111101001001","1110011001010","1111001111010","0000100101101","0000101101100","0000000101000","1111111001100","0000000101101","1111111100110","1111101010010","1111110011000","0000001011101","0000001111101","0000000001111","1111111101100","0000000010010","1111111110101","1111110110101","1111111010011","0000000101001","0000000110111","0000000000111","1111111110111","0000000001000"),
("0000000000111","1111111111000","0000000110110","1111111000100","0000000001100","1111111110011","0000001010010","1111110100101","0000000010001","1111111101101","0000001111100","1111101110111","0000000011010","1111111100011","0000011000000","1111100101000","0000000101010","1111111001111","0000101001110","1111001110000","0000001010101","1111110010010","0001110000110","1101000011010","0001100001011","0001100001011","1101000011010","0001110000110","1111110010010","0000001010101","1111001110000","0000101001110","1111111001111","0000000101010","1111100101000","0000011000000","1111111100011","0000000011010","1111101110111","0000001111100","1111111101101","0000000010001","1111110100101","0000001010010","1111111110011","0000000001100","1111111000100","0000000110110","1111111111000","0000000000111"));


-- components 

-- The samples come from the main main 
-- The Coefficents will be here or in the package 

-- serialfilter component 
COMPONENT serial_filter IS 
  GENERIC(
        NUM_OF_COEFFS : NATURAL );
    PORT( 
        clk     : IN STD_LOGIC;
        reset   : IN STD_LOGIC;
        CO      : IN coefficient_type;
        CE      : IN STD_LOGIC;
        sample1 : IN sample;
        sample2 : IN sample;
        Q	      : OUT Multi_Result);
END COMPONENT;

-- signals 
--SIGNAL CE_FIR1,OE_FIR1,CE_FIR2,OE_FIR2: STD_LOGIC; Not used ?? /shwan
SIGNAL Q_FIR1, Q_FIR2 :  Multi_Result;
SIGNAL CO_FIR1,CO_FIR2 : coefficient_type;

SIGNAL start_filter : STD_LOGIC;

BEGIN 
-- component instantiation 
FIR1:  serial_filter 
    GENERIC MAP (
        NUM_OF_COEFFS => NUM_OF_COEFFS)
    PORT MAP(
        clk => clk,
        reset => updated,
        CO => CO_FIR1,
        CE => start_filter,
        sample1 => sample1,
        sample2 => sample2,
        Q => Q_FIR1);
    
FIR2:  serial_filter
    GENERIC MAP (
        NUM_OF_COEFFS => NUM_OF_COEFFS)
    PORT MAP(
        clk => clk,
        reset => updated,
        CO => CO_FIR2,
        CE => start_filter,
        sample1 => sample1,
        sample2 => sample2,
        Q => Q_FIR2);

PROCESS(clk, updated)
    VARIABLE count : NATURAL RANGE 0 TO NUM_OF_COEFFS;
    VARIABLE count_filters : NATURAL RANGE 0 TO NUM_OF_BANDS+1;
    TYPE state_type IS (IDLE, READ_SAMPLE, UPDATE_FILTER, UPDATE_OUTPUT);
    VARIABLE state : state_type;
    VARIABLE Q_sig : Multi_Result_array;
BEGIN

IF clk'EVENT AND clk = '1' THEN
    IF updated = '1' THEN
        state := READ_SAMPLE;
        count := 0;
        count_filters := 0;
        start_filter <= '0';
        done <= '0';
    ELSE
            CASE (state) IS
                WHEN IDLE =>
                    done <= '0';
                WHEN READ_SAMPLE =>
                    next_sample <= '1';
                    start_filter <= '0';
                    sample_nr <= STD_LOGIC_VECTOR(TO_UNSIGNED(count, 7));
                    state := UPDATE_FILTER;
                    
                WHEN UPDATE_FILTER =>
                    next_sample <= '0';
                    CO_FIR1 <= CO(count_filters, count);
                    CO_FIR2 <= CO(count_filters+1, count);
                    start_filter <= '1';
                    IF count < NUM_OF_COEFFS-1 THEN
                        count := count + 1;
                        state := READ_SAMPLE;
                    ELSE
                        count := 0;
                        state := UPDATE_OUTPUT;
                    END IF;
                    
                WHEN UPDATE_OUTPUT =>
                    Q_sig(count_filters) := Q_FIR1;
                    Q_sig(count_filters+1) := Q_FIR2;
                    start_filter <= '0';
                    IF count_filters < NUM_OF_BANDS-2 THEN
                        count_filters := count_filters + 2; -- since we calculate 2 filters at the time
                        state := READ_SAMPLE;
                    ELSE
                        done <= '1';
                        count_filters := 0;
						Q <= Q_sig;
                        state := IDLE;
                    END IF;
            END CASE;
        END IF;
END IF; --clk
END PROCESS;

END ARCHITECTURE;
