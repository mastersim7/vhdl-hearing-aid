LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.EQ_data_type.all;

ENTITY coeff_io IS
    GENERIC ( 	    N : NATURAL := 24;
		    NUM_OF_TAPS_HALF: NATURAL :=111); -- width of samples and filter coefficients

    PORT (clk     : IN STD_LOGIC;
			 x 	   : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
			 y 	   : IN STD_LOGIC_VECTOR(6 DOWNTO 0); 
			 output  : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)); 
END coeff_io;



ARCHITECTURE coeff_io_arch OF coeff_io IS
TYPE taps_type_2 IS ARRAY(1 TO 2, 1 TO 6) OF STD_LOGIC_VECTOR(23 DOWNTO 0);
CONSTANT tc : taps_type_2 :=
-- Filter coefficients
-- 1
(("111111111111001000011100",
"111111111111000010111011",
"111111111110111101000111",
"111111111110110110111101",
"111111111110110000011001",
"111111111110101001010110"),
-- 2
("111111111111001000011100",
"111111111111000010111011",
"111111111110111101000111",
"111111111110110110111101",
"111111111110110000011001",
"111111111110101001010110"));

BEGIN
	read_coeff: PROCESS(clk, x, y)
	BEGIN
		output <= tc(TO_INTEGER(UNSIGNED(x)),TO_INTEGER(UNSIGNED(y)));
	END PROCESS;
END coeff_io_arch;
