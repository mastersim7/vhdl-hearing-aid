library IEEE;
use IEEE.std_logic_1164.all;

entity sdtb is
end entity;

architecture arch_sdtb of sdtb is

component sd is
  port ( input :in std_logic_vector(11 downto 0); 
         clk :in std_logic; 
         output,add1,add2,latch1 : out std_logic_vector(11 downto 0);
         sign: out std_logic);
end component;

type vals IS ARRAY (0 to 99) of std_logic_vector(11 downto 0); 

constant sin: vals := (
"011111111111",
"100110010100",
"101100011010",
"110010000000",
"110110111000",
"111010110110",
"111101110000",
"111111011111",
"111111111101",
"111111001011",
"111101001010",
"111001111110",
"110101110001",
"110000101100",
"101010111101",
"100100110011",
"011110011100",
"011000001001",
"010010001010",
"001100101110",
"001000000010",
"000100010100",
"000001101100",
"000000010000",
"000000000101",
"000001001011",
"000011011111",
"000110111100",
"001011011000",
"010000101000",
"010110011111",
"011100101110",
"100011000110",
"101001010101",
"101111001101",
"110100011110",
"111000111100",
"111100011010",
"111110110000",
"111111111000",
"111111101111",
"111110010110",
"111011101111",
"111000000010",
"110011011001",
"101101111110",
"100111111111",
"100001101101",
"011011010110",
"010101001010",
"001111011011",
"001010010101",
"000110000110",
"000010111001",
"000000110101",
"000000000001",
"000000011110",
"000010001010",
"000101000010",
"001000111111",
"001101110110",
"010011011011",
"011001011111",
"011111110101",
"100110001010",
"101100010000",
"110001110111",
"110110110001",
"111010110000",
"111101101100",
"111111011101",
"111111111110",
"111111001101",
"111101001110",
"111010000100",
"110101111000",
"110000110101",
"101011000111",
"100100111101",
"011110100110",
"011000010011",
"010010010011",
"001100110110",
"001000001001",
"000100011001",
"000001101111",
"000000010010",
"000000000101",
"000001001001",
"000011011011",
"000110110101",
"001011010000",
"010000011111",
"010110010101",
"011100100100",
"100010111011",
"101001001011",
"101111000100",
"110100010110",
"111000110101"


);





signal input: std_logic_vector(11 downto 0);
signal clk,sign : std_logic:='0'; 
signal output,add1,add2,latch1 : std_logic_vector(11 downto 0);

signal index : integer range 0 to 99:=0;

begin

  clk<= not clk after 100 ns;
  
  S0: SD port map(input, clk, output,add1,add2,latch1, sign);
  
  p0: process
    VARIABLE temp : STD_LOGIC_VECTOR(11 DOWNTO 0);
  begin 

    for i in 0 to 100 loop
      temp := sin(index);
      input <= not temp(12-1) & temp(12-2 downto 0); 
      index<=index+1;
      wait for 1600 ns;
    end loop;
  end process;
end architecture;