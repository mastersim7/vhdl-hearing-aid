library ieee;
use ieee.std_logic_1164.all;

package sine_package is

  constant max_table_value: integer := 2047;
  subtype table_value_type is integer range 0 to max_table_value;

  constant max_table_index: integer := 1023;
  subtype table_index_type is integer range 0 to max_table_index;

  subtype sine_vector_type is std_logic_vector( 11 downto 0 );

  function get_table_value (table_index: table_index_type) return table_value_type;

end;

package body sine_package is

  function get_table_value (table_index: table_index_type) return table_value_type is
    variable table_value: table_value_type;
  begin
    case table_index is
      when 0 =>
        table_value := 2;
      when 1 =>
        table_value := 5;
      when 2 =>
        table_value := 8;
      when 3 =>
        table_value := 11;
      when 4 =>
        table_value := 14;
      when 5 =>
        table_value := 17;
      when 6 =>
        table_value := 20;
      when 7 =>
        table_value := 24;
      when 8 =>
        table_value := 27;
      when 9 =>
        table_value := 30;
      when 10 =>
        table_value := 33;
      when 11 =>
        table_value := 36;
      when 12 =>
        table_value := 39;
      when 13 =>
        table_value := 42;
      when 14 =>
        table_value := 46;
      when 15 =>
        table_value := 49;
      when 16 =>
        table_value := 52;
      when 17 =>
        table_value := 55;
      when 18 =>
        table_value := 58;
      when 19 =>
        table_value := 61;
      when 20 =>
        table_value := 64;
      when 21 =>
        table_value := 67;
      when 22 =>
        table_value := 71;
      when 23 =>
        table_value := 74;
      when 24 =>
        table_value := 77;
      when 25 =>
        table_value := 80;
      when 26 =>
        table_value := 83;
      when 27 =>
        table_value := 86;
      when 28 =>
        table_value := 89;
      when 29 =>
        table_value := 93;
      when 30 =>
        table_value := 96;
      when 31 =>
        table_value := 99;
      when 32 =>
        table_value := 102;
      when 33 =>
        table_value := 105;
      when 34 =>
        table_value := 108;
      when 35 =>
        table_value := 111;
      when 36 =>
        table_value := 115;
      when 37 =>
        table_value := 118;
      when 38 =>
        table_value := 121;
      when 39 =>
        table_value := 124;
      when 40 =>
        table_value := 127;
      when 41 =>
        table_value := 130;
      when 42 =>
        table_value := 133;
      when 43 =>
        table_value := 136;
      when 44 =>
        table_value := 140;
      when 45 =>
        table_value := 143;
      when 46 =>
        table_value := 146;
      when 47 =>
        table_value := 149;
      when 48 =>
        table_value := 152;
      when 49 =>
        table_value := 155;
      when 50 =>
        table_value := 158;
      when 51 =>
        table_value := 162;
      when 52 =>
        table_value := 165;
      when 53 =>
        table_value := 168;
      when 54 =>
        table_value := 171;
      when 55 =>
        table_value := 174;
      when 56 =>
        table_value := 177;
      when 57 =>
        table_value := 180;
      when 58 =>
        table_value := 183;
      when 59 =>
        table_value := 187;
      when 60 =>
        table_value := 190;
      when 61 =>
        table_value := 193;
      when 62 =>
        table_value := 196;
      when 63 =>
        table_value := 199;
      when 64 =>
        table_value := 202;
      when 65 =>
        table_value := 205;
      when 66 =>
        table_value := 208;
      when 67 =>
        table_value := 212;
      when 68 =>
        table_value := 215;
      when 69 =>
        table_value := 218;
      when 70 =>
        table_value := 221;
      when 71 =>
        table_value := 224;
      when 72 =>
        table_value := 227;
      when 73 =>
        table_value := 230;
      when 74 =>
        table_value := 233;
      when 75 =>
        table_value := 237;
      when 76 =>
        table_value := 240;
      when 77 =>
        table_value := 243;
      when 78 =>
        table_value := 246;
      when 79 =>
        table_value := 249;
      when 80 =>
        table_value := 252;
      when 81 =>
        table_value := 255;
      when 82 =>
        table_value := 258;
      when 83 =>
        table_value := 261;
      when 84 =>
        table_value := 265;
      when 85 =>
        table_value := 268;
      when 86 =>
        table_value := 271;
      when 87 =>
        table_value := 274;
      when 88 =>
        table_value := 277;
      when 89 =>
        table_value := 280;
      when 90 =>
        table_value := 283;
      when 91 =>
        table_value := 286;
      when 92 =>
        table_value := 289;
      when 93 =>
        table_value := 293;
      when 94 =>
        table_value := 296;
      when 95 =>
        table_value := 299;
      when 96 =>
        table_value := 302;
      when 97 =>
        table_value := 305;
      when 98 =>
        table_value := 308;
      when 99 =>
        table_value := 311;
      when 100 =>
        table_value := 314;
      when 101 =>
        table_value := 317;
      when 102 =>
        table_value := 321;
      when 103 =>
        table_value := 324;
      when 104 =>
        table_value := 327;
      when 105 =>
        table_value := 330;
      when 106 =>
        table_value := 333;
      when 107 =>
        table_value := 336;
      when 108 =>
        table_value := 339;
      when 109 =>
        table_value := 342;
      when 110 =>
        table_value := 345;
      when 111 =>
        table_value := 348;
      when 112 =>
        table_value := 352;
      when 113 =>
        table_value := 355;
      when 114 =>
        table_value := 358;
      when 115 =>
        table_value := 361;
      when 116 =>
        table_value := 364;
      when 117 =>
        table_value := 367;
      when 118 =>
        table_value := 370;
      when 119 =>
        table_value := 373;
      when 120 =>
        table_value := 376;
      when 121 =>
        table_value := 379;
      when 122 =>
        table_value := 382;
      when 123 =>
        table_value := 385;
      when 124 =>
        table_value := 389;
      when 125 =>
        table_value := 392;
      when 126 =>
        table_value := 395;
      when 127 =>
        table_value := 398;
      when 128 =>
        table_value := 401;
      when 129 =>
        table_value := 404;
      when 130 =>
        table_value := 407;
      when 131 =>
        table_value := 410;
      when 132 =>
        table_value := 413;
      when 133 =>
        table_value := 416;
      when 134 =>
        table_value := 419;
      when 135 =>
        table_value := 422;
      when 136 =>
        table_value := 425;
      when 137 =>
        table_value := 429;
      when 138 =>
        table_value := 432;
      when 139 =>
        table_value := 435;
      when 140 =>
        table_value := 438;
      when 141 =>
        table_value := 441;
      when 142 =>
        table_value := 444;
      when 143 =>
        table_value := 447;
      when 144 =>
        table_value := 450;
      when 145 =>
        table_value := 453;
      when 146 =>
        table_value := 456;
      when 147 =>
        table_value := 459;
      when 148 =>
        table_value := 462;
      when 149 =>
        table_value := 465;
      when 150 =>
        table_value := 468;
      when 151 =>
        table_value := 471;
      when 152 =>
        table_value := 475;
      when 153 =>
        table_value := 478;
      when 154 =>
        table_value := 481;
      when 155 =>
        table_value := 484;
      when 156 =>
        table_value := 487;
      when 157 =>
        table_value := 490;
      when 158 =>
        table_value := 493;
      when 159 =>
        table_value := 496;
      when 160 =>
        table_value := 499;
      when 161 =>
        table_value := 502;
      when 162 =>
        table_value := 505;
      when 163 =>
        table_value := 508;
      when 164 =>
        table_value := 511;
      when 165 =>
        table_value := 514;
      when 166 =>
        table_value := 517;
      when 167 =>
        table_value := 520;
      when 168 =>
        table_value := 523;
      when 169 =>
        table_value := 526;
      when 170 =>
        table_value := 529;
      when 171 =>
        table_value := 532;
      when 172 =>
        table_value := 535;
      when 173 =>
        table_value := 538;
      when 174 =>
        table_value := 541;
      when 175 =>
        table_value := 544;
      when 176 =>
        table_value := 547;
      when 177 =>
        table_value := 550;
      when 178 =>
        table_value := 554;
      when 179 =>
        table_value := 557;
      when 180 =>
        table_value := 560;
      when 181 =>
        table_value := 563;
      when 182 =>
        table_value := 566;
      when 183 =>
        table_value := 569;
      when 184 =>
        table_value := 572;
      when 185 =>
        table_value := 575;
      when 186 =>
        table_value := 578;
      when 187 =>
        table_value := 581;
      when 188 =>
        table_value := 584;
      when 189 =>
        table_value := 587;
      when 190 =>
        table_value := 590;
      when 191 =>
        table_value := 593;
      when 192 =>
        table_value := 596;
      when 193 =>
        table_value := 599;
      when 194 =>
        table_value := 602;
      when 195 =>
        table_value := 605;
      when 196 =>
        table_value := 608;
      when 197 =>
        table_value := 611;
      when 198 =>
        table_value := 614;
      when 199 =>
        table_value := 617;
      when 200 =>
        table_value := 620;
      when 201 =>
        table_value := 623;
      when 202 =>
        table_value := 626;
      when 203 =>
        table_value := 629;
      when 204 =>
        table_value := 632;
      when 205 =>
        table_value := 635;
      when 206 =>
        table_value := 638;
      when 207 =>
        table_value := 641;
      when 208 =>
        table_value := 644;
      when 209 =>
        table_value := 647;
      when 210 =>
        table_value := 650;
      when 211 =>
        table_value := 653;
      when 212 =>
        table_value := 656;
      when 213 =>
        table_value := 658;
      when 214 =>
        table_value := 661;
      when 215 =>
        table_value := 664;
      when 216 =>
        table_value := 667;
      when 217 =>
        table_value := 670;
      when 218 =>
        table_value := 673;
      when 219 =>
        table_value := 676;
      when 220 =>
        table_value := 679;
      when 221 =>
        table_value := 682;
      when 222 =>
        table_value := 685;
      when 223 =>
        table_value := 688;
      when 224 =>
        table_value := 691;
      when 225 =>
        table_value := 694;
      when 226 =>
        table_value := 697;
      when 227 =>
        table_value := 700;
      when 228 =>
        table_value := 703;
      when 229 =>
        table_value := 706;
      when 230 =>
        table_value := 709;
      when 231 =>
        table_value := 712;
      when 232 =>
        table_value := 715;
      when 233 =>
        table_value := 718;
      when 234 =>
        table_value := 721;
      when 235 =>
        table_value := 724;
      when 236 =>
        table_value := 726;
      when 237 =>
        table_value := 729;
      when 238 =>
        table_value := 732;
      when 239 =>
        table_value := 735;
      when 240 =>
        table_value := 738;
      when 241 =>
        table_value := 741;
      when 242 =>
        table_value := 744;
      when 243 =>
        table_value := 747;
      when 244 =>
        table_value := 750;
      when 245 =>
        table_value := 753;
      when 246 =>
        table_value := 756;
      when 247 =>
        table_value := 759;
      when 248 =>
        table_value := 762;
      when 249 =>
        table_value := 764;
      when 250 =>
        table_value := 767;
      when 251 =>
        table_value := 770;
      when 252 =>
        table_value := 773;
      when 253 =>
        table_value := 776;
      when 254 =>
        table_value := 779;
      when 255 =>
        table_value := 782;
      when 256 =>
        table_value := 785;
      when 257 =>
        table_value := 788;
      when 258 =>
        table_value := 791;
      when 259 =>
        table_value := 793;
      when 260 =>
        table_value := 796;
      when 261 =>
        table_value := 799;
      when 262 =>
        table_value := 802;
      when 263 =>
        table_value := 805;
      when 264 =>
        table_value := 808;
      when 265 =>
        table_value := 811;
      when 266 =>
        table_value := 814;
      when 267 =>
        table_value := 817;
      when 268 =>
        table_value := 819;
      when 269 =>
        table_value := 822;
      when 270 =>
        table_value := 825;
      when 271 =>
        table_value := 828;
      when 272 =>
        table_value := 831;
      when 273 =>
        table_value := 834;
      when 274 =>
        table_value := 837;
      when 275 =>
        table_value := 840;
      when 276 =>
        table_value := 842;
      when 277 =>
        table_value := 845;
      when 278 =>
        table_value := 848;
      when 279 =>
        table_value := 851;
      when 280 =>
        table_value := 854;
      when 281 =>
        table_value := 857;
      when 282 =>
        table_value := 860;
      when 283 =>
        table_value := 862;
      when 284 =>
        table_value := 865;
      when 285 =>
        table_value := 868;
      when 286 =>
        table_value := 871;
      when 287 =>
        table_value := 874;
      when 288 =>
        table_value := 877;
      when 289 =>
        table_value := 879;
      when 290 =>
        table_value := 882;
      when 291 =>
        table_value := 885;
      when 292 =>
        table_value := 888;
      when 293 =>
        table_value := 891;
      when 294 =>
        table_value := 894;
      when 295 =>
        table_value := 896;
      when 296 =>
        table_value := 899;
      when 297 =>
        table_value := 902;
      when 298 =>
        table_value := 905;
      when 299 =>
        table_value := 908;
      when 300 =>
        table_value := 911;
      when 301 =>
        table_value := 913;
      when 302 =>
        table_value := 916;
      when 303 =>
        table_value := 919;
      when 304 =>
        table_value := 922;
      when 305 =>
        table_value := 925;
      when 306 =>
        table_value := 927;
      when 307 =>
        table_value := 930;
      when 308 =>
        table_value := 933;
      when 309 =>
        table_value := 936;
      when 310 =>
        table_value := 939;
      when 311 =>
        table_value := 941;
      when 312 =>
        table_value := 944;
      when 313 =>
        table_value := 947;
      when 314 =>
        table_value := 950;
      when 315 =>
        table_value := 952;
      when 316 =>
        table_value := 955;
      when 317 =>
        table_value := 958;
      when 318 =>
        table_value := 961;
      when 319 =>
        table_value := 964;
      when 320 =>
        table_value := 966;
      when 321 =>
        table_value := 969;
      when 322 =>
        table_value := 972;
      when 323 =>
        table_value := 975;
      when 324 =>
        table_value := 977;
      when 325 =>
        table_value := 980;
      when 326 =>
        table_value := 983;
      when 327 =>
        table_value := 986;
      when 328 =>
        table_value := 988;
      when 329 =>
        table_value := 991;
      when 330 =>
        table_value := 994;
      when 331 =>
        table_value := 997;
      when 332 =>
        table_value := 999;
      when 333 =>
        table_value := 1002;
      when 334 =>
        table_value := 1005;
      when 335 =>
        table_value := 1008;
      when 336 =>
        table_value := 1010;
      when 337 =>
        table_value := 1013;
      when 338 =>
        table_value := 1016;
      when 339 =>
        table_value := 1019;
      when 340 =>
        table_value := 1021;
      when 341 =>
        table_value := 1024;
      when 342 =>
        table_value := 1027;
      when 343 =>
        table_value := 1029;
      when 344 =>
        table_value := 1032;
      when 345 =>
        table_value := 1035;
      when 346 =>
        table_value := 1038;
      when 347 =>
        table_value := 1040;
      when 348 =>
        table_value := 1043;
      when 349 =>
        table_value := 1046;
      when 350 =>
        table_value := 1048;
      when 351 =>
        table_value := 1051;
      when 352 =>
        table_value := 1054;
      when 353 =>
        table_value := 1056;
      when 354 =>
        table_value := 1059;
      when 355 =>
        table_value := 1062;
      when 356 =>
        table_value := 1064;
      when 357 =>
        table_value := 1067;
      when 358 =>
        table_value := 1070;
      when 359 =>
        table_value := 1072;
      when 360 =>
        table_value := 1075;
      when 361 =>
        table_value := 1078;
      when 362 =>
        table_value := 1081;
      when 363 =>
        table_value := 1083;
      when 364 =>
        table_value := 1086;
      when 365 =>
        table_value := 1088;
      when 366 =>
        table_value := 1091;
      when 367 =>
        table_value := 1094;
      when 368 =>
        table_value := 1096;
      when 369 =>
        table_value := 1099;
      when 370 =>
        table_value := 1102;
      when 371 =>
        table_value := 1104;
      when 372 =>
        table_value := 1107;
      when 373 =>
        table_value := 1110;
      when 374 =>
        table_value := 1112;
      when 375 =>
        table_value := 1115;
      when 376 =>
        table_value := 1118;
      when 377 =>
        table_value := 1120;
      when 378 =>
        table_value := 1123;
      when 379 =>
        table_value := 1125;
      when 380 =>
        table_value := 1128;
      when 381 =>
        table_value := 1131;
      when 382 =>
        table_value := 1133;
      when 383 =>
        table_value := 1136;
      when 384 =>
        table_value := 1139;
      when 385 =>
        table_value := 1141;
      when 386 =>
        table_value := 1144;
      when 387 =>
        table_value := 1146;
      when 388 =>
        table_value := 1149;
      when 389 =>
        table_value := 1152;
      when 390 =>
        table_value := 1154;
      when 391 =>
        table_value := 1157;
      when 392 =>
        table_value := 1159;
      when 393 =>
        table_value := 1162;
      when 394 =>
        table_value := 1165;
      when 395 =>
        table_value := 1167;
      when 396 =>
        table_value := 1170;
      when 397 =>
        table_value := 1172;
      when 398 =>
        table_value := 1175;
      when 399 =>
        table_value := 1177;
      when 400 =>
        table_value := 1180;
      when 401 =>
        table_value := 1183;
      when 402 =>
        table_value := 1185;
      when 403 =>
        table_value := 1188;
      when 404 =>
        table_value := 1190;
      when 405 =>
        table_value := 1193;
      when 406 =>
        table_value := 1195;
      when 407 =>
        table_value := 1198;
      when 408 =>
        table_value := 1200;
      when 409 =>
        table_value := 1203;
      when 410 =>
        table_value := 1205;
      when 411 =>
        table_value := 1208;
      when 412 =>
        table_value := 1211;
      when 413 =>
        table_value := 1213;
      when 414 =>
        table_value := 1216;
      when 415 =>
        table_value := 1218;
      when 416 =>
        table_value := 1221;
      when 417 =>
        table_value := 1223;
      when 418 =>
        table_value := 1226;
      when 419 =>
        table_value := 1228;
      when 420 =>
        table_value := 1231;
      when 421 =>
        table_value := 1233;
      when 422 =>
        table_value := 1236;
      when 423 =>
        table_value := 1238;
      when 424 =>
        table_value := 1241;
      when 425 =>
        table_value := 1243;
      when 426 =>
        table_value := 1246;
      when 427 =>
        table_value := 1248;
      when 428 =>
        table_value := 1251;
      when 429 =>
        table_value := 1253;
      when 430 =>
        table_value := 1256;
      when 431 =>
        table_value := 1258;
      when 432 =>
        table_value := 1261;
      when 433 =>
        table_value := 1263;
      when 434 =>
        table_value := 1266;
      when 435 =>
        table_value := 1268;
      when 436 =>
        table_value := 1270;
      when 437 =>
        table_value := 1273;
      when 438 =>
        table_value := 1275;
      when 439 =>
        table_value := 1278;
      when 440 =>
        table_value := 1280;
      when 441 =>
        table_value := 1283;
      when 442 =>
        table_value := 1285;
      when 443 =>
        table_value := 1288;
      when 444 =>
        table_value := 1290;
      when 445 =>
        table_value := 1293;
      when 446 =>
        table_value := 1295;
      when 447 =>
        table_value := 1297;
      when 448 =>
        table_value := 1300;
      when 449 =>
        table_value := 1302;
      when 450 =>
        table_value := 1305;
      when 451 =>
        table_value := 1307;
      when 452 =>
        table_value := 1309;
      when 453 =>
        table_value := 1312;
      when 454 =>
        table_value := 1314;
      when 455 =>
        table_value := 1317;
      when 456 =>
        table_value := 1319;
      when 457 =>
        table_value := 1322;
      when 458 =>
        table_value := 1324;
      when 459 =>
        table_value := 1326;
      when 460 =>
        table_value := 1329;
      when 461 =>
        table_value := 1331;
      when 462 =>
        table_value := 1333;
      when 463 =>
        table_value := 1336;
      when 464 =>
        table_value := 1338;
      when 465 =>
        table_value := 1341;
      when 466 =>
        table_value := 1343;
      when 467 =>
        table_value := 1345;
      when 468 =>
        table_value := 1348;
      when 469 =>
        table_value := 1350;
      when 470 =>
        table_value := 1352;
      when 471 =>
        table_value := 1355;
      when 472 =>
        table_value := 1357;
      when 473 =>
        table_value := 1359;
      when 474 =>
        table_value := 1362;
      when 475 =>
        table_value := 1364;
      when 476 =>
        table_value := 1367;
      when 477 =>
        table_value := 1369;
      when 478 =>
        table_value := 1371;
      when 479 =>
        table_value := 1374;
      when 480 =>
        table_value := 1376;
      when 481 =>
        table_value := 1378;
      when 482 =>
        table_value := 1380;
      when 483 =>
        table_value := 1383;
      when 484 =>
        table_value := 1385;
      when 485 =>
        table_value := 1387;
      when 486 =>
        table_value := 1390;
      when 487 =>
        table_value := 1392;
      when 488 =>
        table_value := 1394;
      when 489 =>
        table_value := 1397;
      when 490 =>
        table_value := 1399;
      when 491 =>
        table_value := 1401;
      when 492 =>
        table_value := 1404;
      when 493 =>
        table_value := 1406;
      when 494 =>
        table_value := 1408;
      when 495 =>
        table_value := 1410;
      when 496 =>
        table_value := 1413;
      when 497 =>
        table_value := 1415;
      when 498 =>
        table_value := 1417;
      when 499 =>
        table_value := 1419;
      when 500 =>
        table_value := 1422;
      when 501 =>
        table_value := 1424;
      when 502 =>
        table_value := 1426;
      when 503 =>
        table_value := 1428;
      when 504 =>
        table_value := 1431;
      when 505 =>
        table_value := 1433;
      when 506 =>
        table_value := 1435;
      when 507 =>
        table_value := 1437;
      when 508 =>
        table_value := 1440;
      when 509 =>
        table_value := 1442;
      when 510 =>
        table_value := 1444;
      when 511 =>
        table_value := 1446;
      when 512 =>
        table_value := 1449;
      when 513 =>
        table_value := 1451;
      when 514 =>
        table_value := 1453;
      when 515 =>
        table_value := 1455;
      when 516 =>
        table_value := 1457;
      when 517 =>
        table_value := 1460;
      when 518 =>
        table_value := 1462;
      when 519 =>
        table_value := 1464;
      when 520 =>
        table_value := 1466;
      when 521 =>
        table_value := 1468;
      when 522 =>
        table_value := 1471;
      when 523 =>
        table_value := 1473;
      when 524 =>
        table_value := 1475;
      when 525 =>
        table_value := 1477;
      when 526 =>
        table_value := 1479;
      when 527 =>
        table_value := 1481;
      when 528 =>
        table_value := 1484;
      when 529 =>
        table_value := 1486;
      when 530 =>
        table_value := 1488;
      when 531 =>
        table_value := 1490;
      when 532 =>
        table_value := 1492;
      when 533 =>
        table_value := 1494;
      when 534 =>
        table_value := 1497;
      when 535 =>
        table_value := 1499;
      when 536 =>
        table_value := 1501;
      when 537 =>
        table_value := 1503;
      when 538 =>
        table_value := 1505;
      when 539 =>
        table_value := 1507;
      when 540 =>
        table_value := 1509;
      when 541 =>
        table_value := 1511;
      when 542 =>
        table_value := 1514;
      when 543 =>
        table_value := 1516;
      when 544 =>
        table_value := 1518;
      when 545 =>
        table_value := 1520;
      when 546 =>
        table_value := 1522;
      when 547 =>
        table_value := 1524;
      when 548 =>
        table_value := 1526;
      when 549 =>
        table_value := 1528;
      when 550 =>
        table_value := 1530;
      when 551 =>
        table_value := 1532;
      when 552 =>
        table_value := 1535;
      when 553 =>
        table_value := 1537;
      when 554 =>
        table_value := 1539;
      when 555 =>
        table_value := 1541;
      when 556 =>
        table_value := 1543;
      when 557 =>
        table_value := 1545;
      when 558 =>
        table_value := 1547;
      when 559 =>
        table_value := 1549;
      when 560 =>
        table_value := 1551;
      when 561 =>
        table_value := 1553;
      when 562 =>
        table_value := 1555;
      when 563 =>
        table_value := 1557;
      when 564 =>
        table_value := 1559;
      when 565 =>
        table_value := 1561;
      when 566 =>
        table_value := 1563;
      when 567 =>
        table_value := 1565;
      when 568 =>
        table_value := 1567;
      when 569 =>
        table_value := 1569;
      when 570 =>
        table_value := 1571;
      when 571 =>
        table_value := 1573;
      when 572 =>
        table_value := 1575;
      when 573 =>
        table_value := 1577;
      when 574 =>
        table_value := 1579;
      when 575 =>
        table_value := 1581;
      when 576 =>
        table_value := 1583;
      when 577 =>
        table_value := 1585;
      when 578 =>
        table_value := 1587;
      when 579 =>
        table_value := 1589;
      when 580 =>
        table_value := 1591;
      when 581 =>
        table_value := 1593;
      when 582 =>
        table_value := 1595;
      when 583 =>
        table_value := 1597;
      when 584 =>
        table_value := 1599;
      when 585 =>
        table_value := 1601;
      when 586 =>
        table_value := 1603;
      when 587 =>
        table_value := 1605;
      when 588 =>
        table_value := 1607;
      when 589 =>
        table_value := 1609;
      when 590 =>
        table_value := 1611;
      when 591 =>
        table_value := 1613;
      when 592 =>
        table_value := 1615;
      when 593 =>
        table_value := 1617;
      when 594 =>
        table_value := 1619;
      when 595 =>
        table_value := 1620;
      when 596 =>
        table_value := 1622;
      when 597 =>
        table_value := 1624;
      when 598 =>
        table_value := 1626;
      when 599 =>
        table_value := 1628;
      when 600 =>
        table_value := 1630;
      when 601 =>
        table_value := 1632;
      when 602 =>
        table_value := 1634;
      when 603 =>
        table_value := 1636;
      when 604 =>
        table_value := 1638;
      when 605 =>
        table_value := 1639;
      when 606 =>
        table_value := 1641;
      when 607 =>
        table_value := 1643;
      when 608 =>
        table_value := 1645;
      when 609 =>
        table_value := 1647;
      when 610 =>
        table_value := 1649;
      when 611 =>
        table_value := 1651;
      when 612 =>
        table_value := 1653;
      when 613 =>
        table_value := 1654;
      when 614 =>
        table_value := 1656;
      when 615 =>
        table_value := 1658;
      when 616 =>
        table_value := 1660;
      when 617 =>
        table_value := 1662;
      when 618 =>
        table_value := 1664;
      when 619 =>
        table_value := 1665;
      when 620 =>
        table_value := 1667;
      when 621 =>
        table_value := 1669;
      when 622 =>
        table_value := 1671;
      when 623 =>
        table_value := 1673;
      when 624 =>
        table_value := 1674;
      when 625 =>
        table_value := 1676;
      when 626 =>
        table_value := 1678;
      when 627 =>
        table_value := 1680;
      when 628 =>
        table_value := 1682;
      when 629 =>
        table_value := 1683;
      when 630 =>
        table_value := 1685;
      when 631 =>
        table_value := 1687;
      when 632 =>
        table_value := 1689;
      when 633 =>
        table_value := 1691;
      when 634 =>
        table_value := 1692;
      when 635 =>
        table_value := 1694;
      when 636 =>
        table_value := 1696;
      when 637 =>
        table_value := 1698;
      when 638 =>
        table_value := 1699;
      when 639 =>
        table_value := 1701;
      when 640 =>
        table_value := 1703;
      when 641 =>
        table_value := 1705;
      when 642 =>
        table_value := 1706;
      when 643 =>
        table_value := 1708;
      when 644 =>
        table_value := 1710;
      when 645 =>
        table_value := 1712;
      when 646 =>
        table_value := 1713;
      when 647 =>
        table_value := 1715;
      when 648 =>
        table_value := 1717;
      when 649 =>
        table_value := 1718;
      when 650 =>
        table_value := 1720;
      when 651 =>
        table_value := 1722;
      when 652 =>
        table_value := 1724;
      when 653 =>
        table_value := 1725;
      when 654 =>
        table_value := 1727;
      when 655 =>
        table_value := 1729;
      when 656 =>
        table_value := 1730;
      when 657 =>
        table_value := 1732;
      when 658 =>
        table_value := 1734;
      when 659 =>
        table_value := 1735;
      when 660 =>
        table_value := 1737;
      when 661 =>
        table_value := 1739;
      when 662 =>
        table_value := 1740;
      when 663 =>
        table_value := 1742;
      when 664 =>
        table_value := 1744;
      when 665 =>
        table_value := 1745;
      when 666 =>
        table_value := 1747;
      when 667 =>
        table_value := 1748;
      when 668 =>
        table_value := 1750;
      when 669 =>
        table_value := 1752;
      when 670 =>
        table_value := 1753;
      when 671 =>
        table_value := 1755;
      when 672 =>
        table_value := 1757;
      when 673 =>
        table_value := 1758;
      when 674 =>
        table_value := 1760;
      when 675 =>
        table_value := 1761;
      when 676 =>
        table_value := 1763;
      when 677 =>
        table_value := 1765;
      when 678 =>
        table_value := 1766;
      when 679 =>
        table_value := 1768;
      when 680 =>
        table_value := 1769;
      when 681 =>
        table_value := 1771;
      when 682 =>
        table_value := 1772;
      when 683 =>
        table_value := 1774;
      when 684 =>
        table_value := 1776;
      when 685 =>
        table_value := 1777;
      when 686 =>
        table_value := 1779;
      when 687 =>
        table_value := 1780;
      when 688 =>
        table_value := 1782;
      when 689 =>
        table_value := 1783;
      when 690 =>
        table_value := 1785;
      when 691 =>
        table_value := 1786;
      when 692 =>
        table_value := 1788;
      when 693 =>
        table_value := 1790;
      when 694 =>
        table_value := 1791;
      when 695 =>
        table_value := 1793;
      when 696 =>
        table_value := 1794;
      when 697 =>
        table_value := 1796;
      when 698 =>
        table_value := 1797;
      when 699 =>
        table_value := 1799;
      when 700 =>
        table_value := 1800;
      when 701 =>
        table_value := 1802;
      when 702 =>
        table_value := 1803;
      when 703 =>
        table_value := 1805;
      when 704 =>
        table_value := 1806;
      when 705 =>
        table_value := 1808;
      when 706 =>
        table_value := 1809;
      when 707 =>
        table_value := 1810;
      when 708 =>
        table_value := 1812;
      when 709 =>
        table_value := 1813;
      when 710 =>
        table_value := 1815;
      when 711 =>
        table_value := 1816;
      when 712 =>
        table_value := 1818;
      when 713 =>
        table_value := 1819;
      when 714 =>
        table_value := 1821;
      when 715 =>
        table_value := 1822;
      when 716 =>
        table_value := 1823;
      when 717 =>
        table_value := 1825;
      when 718 =>
        table_value := 1826;
      when 719 =>
        table_value := 1828;
      when 720 =>
        table_value := 1829;
      when 721 =>
        table_value := 1831;
      when 722 =>
        table_value := 1832;
      when 723 =>
        table_value := 1833;
      when 724 =>
        table_value := 1835;
      when 725 =>
        table_value := 1836;
      when 726 =>
        table_value := 1838;
      when 727 =>
        table_value := 1839;
      when 728 =>
        table_value := 1840;
      when 729 =>
        table_value := 1842;
      when 730 =>
        table_value := 1843;
      when 731 =>
        table_value := 1844;
      when 732 =>
        table_value := 1846;
      when 733 =>
        table_value := 1847;
      when 734 =>
        table_value := 1848;
      when 735 =>
        table_value := 1850;
      when 736 =>
        table_value := 1851;
      when 737 =>
        table_value := 1852;
      when 738 =>
        table_value := 1854;
      when 739 =>
        table_value := 1855;
      when 740 =>
        table_value := 1856;
      when 741 =>
        table_value := 1858;
      when 742 =>
        table_value := 1859;
      when 743 =>
        table_value := 1860;
      when 744 =>
        table_value := 1862;
      when 745 =>
        table_value := 1863;
      when 746 =>
        table_value := 1864;
      when 747 =>
        table_value := 1866;
      when 748 =>
        table_value := 1867;
      when 749 =>
        table_value := 1868;
      when 750 =>
        table_value := 1869;
      when 751 =>
        table_value := 1871;
      when 752 =>
        table_value := 1872;
      when 753 =>
        table_value := 1873;
      when 754 =>
        table_value := 1875;
      when 755 =>
        table_value := 1876;
      when 756 =>
        table_value := 1877;
      when 757 =>
        table_value := 1878;
      when 758 =>
        table_value := 1880;
      when 759 =>
        table_value := 1881;
      when 760 =>
        table_value := 1882;
      when 761 =>
        table_value := 1883;
      when 762 =>
        table_value := 1885;
      when 763 =>
        table_value := 1886;
      when 764 =>
        table_value := 1887;
      when 765 =>
        table_value := 1888;
      when 766 =>
        table_value := 1889;
      when 767 =>
        table_value := 1891;
      when 768 =>
        table_value := 1892;
      when 769 =>
        table_value := 1893;
      when 770 =>
        table_value := 1894;
      when 771 =>
        table_value := 1895;
      when 772 =>
        table_value := 1897;
      when 773 =>
        table_value := 1898;
      when 774 =>
        table_value := 1899;
      when 775 =>
        table_value := 1900;
      when 776 =>
        table_value := 1901;
      when 777 =>
        table_value := 1902;
      when 778 =>
        table_value := 1904;
      when 779 =>
        table_value := 1905;
      when 780 =>
        table_value := 1906;
      when 781 =>
        table_value := 1907;
      when 782 =>
        table_value := 1908;
      when 783 =>
        table_value := 1909;
      when 784 =>
        table_value := 1910;
      when 785 =>
        table_value := 1912;
      when 786 =>
        table_value := 1913;
      when 787 =>
        table_value := 1914;
      when 788 =>
        table_value := 1915;
      when 789 =>
        table_value := 1916;
      when 790 =>
        table_value := 1917;
      when 791 =>
        table_value := 1918;
      when 792 =>
        table_value := 1919;
      when 793 =>
        table_value := 1920;
      when 794 =>
        table_value := 1921;
      when 795 =>
        table_value := 1923;
      when 796 =>
        table_value := 1924;
      when 797 =>
        table_value := 1925;
      when 798 =>
        table_value := 1926;
      when 799 =>
        table_value := 1927;
      when 800 =>
        table_value := 1928;
      when 801 =>
        table_value := 1929;
      when 802 =>
        table_value := 1930;
      when 803 =>
        table_value := 1931;
      when 804 =>
        table_value := 1932;
      when 805 =>
        table_value := 1933;
      when 806 =>
        table_value := 1934;
      when 807 =>
        table_value := 1935;
      when 808 =>
        table_value := 1936;
      when 809 =>
        table_value := 1937;
      when 810 =>
        table_value := 1938;
      when 811 =>
        table_value := 1939;
      when 812 =>
        table_value := 1940;
      when 813 =>
        table_value := 1941;
      when 814 =>
        table_value := 1942;
      when 815 =>
        table_value := 1943;
      when 816 =>
        table_value := 1944;
      when 817 =>
        table_value := 1945;
      when 818 =>
        table_value := 1946;
      when 819 =>
        table_value := 1947;
      when 820 =>
        table_value := 1948;
      when 821 =>
        table_value := 1949;
      when 822 =>
        table_value := 1950;
      when 823 =>
        table_value := 1951;
      when 824 =>
        table_value := 1952;
      when 825 =>
        table_value := 1953;
      when 826 =>
        table_value := 1954;
      when 827 =>
        table_value := 1955;
      when 828 =>
        table_value := 1956;
      when 829 =>
        table_value := 1957;
      when 830 =>
        table_value := 1957;
      when 831 =>
        table_value := 1958;
      when 832 =>
        table_value := 1959;
      when 833 =>
        table_value := 1960;
      when 834 =>
        table_value := 1961;
      when 835 =>
        table_value := 1962;
      when 836 =>
        table_value := 1963;
      when 837 =>
        table_value := 1964;
      when 838 =>
        table_value := 1965;
      when 839 =>
        table_value := 1966;
      when 840 =>
        table_value := 1966;
      when 841 =>
        table_value := 1967;
      when 842 =>
        table_value := 1968;
      when 843 =>
        table_value := 1969;
      when 844 =>
        table_value := 1970;
      when 845 =>
        table_value := 1971;
      when 846 =>
        table_value := 1972;
      when 847 =>
        table_value := 1972;
      when 848 =>
        table_value := 1973;
      when 849 =>
        table_value := 1974;
      when 850 =>
        table_value := 1975;
      when 851 =>
        table_value := 1976;
      when 852 =>
        table_value := 1977;
      when 853 =>
        table_value := 1977;
      when 854 =>
        table_value := 1978;
      when 855 =>
        table_value := 1979;
      when 856 =>
        table_value := 1980;
      when 857 =>
        table_value := 1981;
      when 858 =>
        table_value := 1981;
      when 859 =>
        table_value := 1982;
      when 860 =>
        table_value := 1983;
      when 861 =>
        table_value := 1984;
      when 862 =>
        table_value := 1985;
      when 863 =>
        table_value := 1985;
      when 864 =>
        table_value := 1986;
      when 865 =>
        table_value := 1987;
      when 866 =>
        table_value := 1988;
      when 867 =>
        table_value := 1988;
      when 868 =>
        table_value := 1989;
      when 869 =>
        table_value := 1990;
      when 870 =>
        table_value := 1991;
      when 871 =>
        table_value := 1991;
      when 872 =>
        table_value := 1992;
      when 873 =>
        table_value := 1993;
      when 874 =>
        table_value := 1993;
      when 875 =>
        table_value := 1994;
      when 876 =>
        table_value := 1995;
      when 877 =>
        table_value := 1996;
      when 878 =>
        table_value := 1996;
      when 879 =>
        table_value := 1997;
      when 880 =>
        table_value := 1998;
      when 881 =>
        table_value := 1998;
      when 882 =>
        table_value := 1999;
      when 883 =>
        table_value := 2000;
      when 884 =>
        table_value := 2000;
      when 885 =>
        table_value := 2001;
      when 886 =>
        table_value := 2002;
      when 887 =>
        table_value := 2002;
      when 888 =>
        table_value := 2003;
      when 889 =>
        table_value := 2004;
      when 890 =>
        table_value := 2004;
      when 891 =>
        table_value := 2005;
      when 892 =>
        table_value := 2005;
      when 893 =>
        table_value := 2006;
      when 894 =>
        table_value := 2007;
      when 895 =>
        table_value := 2007;
      when 896 =>
        table_value := 2008;
      when 897 =>
        table_value := 2009;
      when 898 =>
        table_value := 2009;
      when 899 =>
        table_value := 2010;
      when 900 =>
        table_value := 2010;
      when 901 =>
        table_value := 2011;
      when 902 =>
        table_value := 2012;
      when 903 =>
        table_value := 2012;
      when 904 =>
        table_value := 2013;
      when 905 =>
        table_value := 2013;
      when 906 =>
        table_value := 2014;
      when 907 =>
        table_value := 2014;
      when 908 =>
        table_value := 2015;
      when 909 =>
        table_value := 2016;
      when 910 =>
        table_value := 2016;
      when 911 =>
        table_value := 2017;
      when 912 =>
        table_value := 2017;
      when 913 =>
        table_value := 2018;
      when 914 =>
        table_value := 2018;
      when 915 =>
        table_value := 2019;
      when 916 =>
        table_value := 2019;
      when 917 =>
        table_value := 2020;
      when 918 =>
        table_value := 2020;
      when 919 =>
        table_value := 2021;
      when 920 =>
        table_value := 2021;
      when 921 =>
        table_value := 2022;
      when 922 =>
        table_value := 2022;
      when 923 =>
        table_value := 2023;
      when 924 =>
        table_value := 2023;
      when 925 =>
        table_value := 2024;
      when 926 =>
        table_value := 2024;
      when 927 =>
        table_value := 2025;
      when 928 =>
        table_value := 2025;
      when 929 =>
        table_value := 2026;
      when 930 =>
        table_value := 2026;
      when 931 =>
        table_value := 2026;
      when 932 =>
        table_value := 2027;
      when 933 =>
        table_value := 2027;
      when 934 =>
        table_value := 2028;
      when 935 =>
        table_value := 2028;
      when 936 =>
        table_value := 2029;
      when 937 =>
        table_value := 2029;
      when 938 =>
        table_value := 2029;
      when 939 =>
        table_value := 2030;
      when 940 =>
        table_value := 2030;
      when 941 =>
        table_value := 2031;
      when 942 =>
        table_value := 2031;
      when 943 =>
        table_value := 2031;
      when 944 =>
        table_value := 2032;
      when 945 =>
        table_value := 2032;
      when 946 =>
        table_value := 2033;
      when 947 =>
        table_value := 2033;
      when 948 =>
        table_value := 2033;
      when 949 =>
        table_value := 2034;
      when 950 =>
        table_value := 2034;
      when 951 =>
        table_value := 2034;
      when 952 =>
        table_value := 2035;
      when 953 =>
        table_value := 2035;
      when 954 =>
        table_value := 2035;
      when 955 =>
        table_value := 2036;
      when 956 =>
        table_value := 2036;
      when 957 =>
        table_value := 2036;
      when 958 =>
        table_value := 2037;
      when 959 =>
        table_value := 2037;
      when 960 =>
        table_value := 2037;
      when 961 =>
        table_value := 2038;
      when 962 =>
        table_value := 2038;
      when 963 =>
        table_value := 2038;
      when 964 =>
        table_value := 2038;
      when 965 =>
        table_value := 2039;
      when 966 =>
        table_value := 2039;
      when 967 =>
        table_value := 2039;
      when 968 =>
        table_value := 2040;
      when 969 =>
        table_value := 2040;
      when 970 =>
        table_value := 2040;
      when 971 =>
        table_value := 2040;
      when 972 =>
        table_value := 2041;
      when 973 =>
        table_value := 2041;
      when 974 =>
        table_value := 2041;
      when 975 =>
        table_value := 2041;
      when 976 =>
        table_value := 2042;
      when 977 =>
        table_value := 2042;
      when 978 =>
        table_value := 2042;
      when 979 =>
        table_value := 2042;
      when 980 =>
        table_value := 2042;
      when 981 =>
        table_value := 2043;
      when 982 =>
        table_value := 2043;
      when 983 =>
        table_value := 2043;
      when 984 =>
        table_value := 2043;
      when 985 =>
        table_value := 2043;
      when 986 =>
        table_value := 2044;
      when 987 =>
        table_value := 2044;
      when 988 =>
        table_value := 2044;
      when 989 =>
        table_value := 2044;
      when 990 =>
        table_value := 2044;
      when 991 =>
        table_value := 2044;
      when 992 =>
        table_value := 2045;
      when 993 =>
        table_value := 2045;
      when 994 =>
        table_value := 2045;
      when 995 =>
        table_value := 2045;
      when 996 =>
        table_value := 2045;
      when 997 =>
        table_value := 2045;
      when 998 =>
        table_value := 2045;
      when 999 =>
        table_value := 2046;
      when 1000 =>
        table_value := 2046;
      when 1001 =>
        table_value := 2046;
      when 1002 =>
        table_value := 2046;
      when 1003 =>
        table_value := 2046;
      when 1004 =>
        table_value := 2046;
      when 1005 =>
        table_value := 2046;
      when 1006 =>
        table_value := 2046;
      when 1007 =>
        table_value := 2046;
      when 1008 =>
        table_value := 2046;
      when 1009 =>
        table_value := 2046;
      when 1010 =>
        table_value := 2047;
      when 1011 =>
        table_value := 2047;
      when 1012 =>
        table_value := 2047;
      when 1013 =>
        table_value := 2047;
      when 1014 =>
        table_value := 2047;
      when 1015 =>
        table_value := 2047;
      when 1016 =>
        table_value := 2047;
      when 1017 =>
        table_value := 2047;
      when 1018 =>
        table_value := 2047;
      when 1019 =>
        table_value := 2047;
      when 1020 =>
        table_value := 2047;
      when 1021 =>
        table_value := 2047;
      when 1022 =>
        table_value := 2047;
      when 1023 =>
        table_value := 2047;
    end case;
    return table_value;
  end;

end;
