-- Description:
-- filterblock_main.vhd
-- Author: Shwan Ciyako,Anandhavel Sakthivel
-- It is still in the implementation phase. 
-- This files adds needed components together to make a filterbank, you are welcome to make changes but make shure to update the whole chain of files that will be affected

-- 2011-03-30, Mathias Lundell
-- Works essentially in the same way. There is still a simulation error which
-- I believe is constrained to simulation and not implementation on fpga.
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_signed.ALL;
USE work.EQ_data_type.ALL;

ENTITY filterblock_main IS
	  GENERIC(
            NUM_BITS_OUT : NATURAL ;
            NUM_OF_SAMPLES : NATURAL ;
            NUM_OF_COEFFS : NATURAL ;
            NUM_OF_BANDS: NATURAL );
    PORT( 
            clk     : IN STD_LOGIC;
            sample1 : IN sample;            
            sample2 : IN sample;
            updated : IN STD_LOGIC; 
            Q       : OUT Multi_Result_array;
            done    : OUT STD_LOGIC;
            next_sample : OUT STD_LOGIC;
            sample_nr : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END filterblock_main;

ARCHITECTURE  filterblock_main_arch OF filterblock_main IS 
-- constants 
CONSTANT CO:taps_type:=
(("0000000010100","0000000010101","0000000010110","0000000010111","0000000011000","0000000011001","0000000011010","0000000011011","0000000011100","0000000011101","0000000011110","0000000011110","0000000011111","0000000100000","0000000100001","0000000100010","0000000100011","0000000100100","0000000100101","0000000100110","0000000100111","0000000101000","0000000101001","0000000101010","0000000101011","0000000101011","0000000101100","0000000101101","0000000101110","0000000101111","0000000101111","0000000110000","0000000110001","0000000110001","0000000110010","0000000110010","0000000110011","0000000110011","0000000110100","0000000110100","0000000110101","0000000110101","0000000110101","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110110","0000000110101","0000000110101","0000000110101","0000000110100","0000000110100","0000000110011","0000000110011","0000000110010","0000000110010","0000000110001","0000000110001","0000000110000","0000000101111","0000000101111","0000000101110","0000000101101","0000000101100","0000000101011","0000000101011","0000000101010","0000000101001","0000000101000","0000000100111","0000000100110","0000000100101","0000000100100","0000000100011","0000000100010","0000000100001","0000000100000","0000000011111","0000000011110","0000000011110","0000000011101","0000000011100","0000000011011","0000000011010","0000000011001","0000000011000","0000000010111","0000000010110","0000000010101","0000000010100"),
("1111111110101","1111111110110","1111111110111","1111111111001","1111111111011","1111111111100","1111111111110","0000000000000","0000000000011","0000000000101","0000000000111","0000000001010","0000000001100","0000000001111","0000000010010","0000000010101","0000000011000","0000000011011","0000000011110","0000000100001","0000000100101","0000000101000","0000000101011","0000000101110","0000000110010","0000000110101","0000000111000","0000000111011","0000000111111","0000001000010","0000001000101","0000001001000","0000001001011","0000001001110","0000001010000","0000001010011","0000001010101","0000001011000","0000001011010","0000001011100","0000001011110","0000001011111","0000001100001","0000001100010","0000001100011","0000001100100","0000001100101","0000001100110","0000001100110","0000001100110","0000001100110","0000001100110","0000001100110","0000001100101","0000001100100","0000001100011","0000001100010","0000001100001","0000001011111","0000001011110","0000001011100","0000001011010","0000001011000","0000001010101","0000001010011","0000001010000","0000001001110","0000001001011","0000001001000","0000001000101","0000001000010","0000000111111","0000000111011","0000000111000","0000000110101","0000000110010","0000000101110","0000000101011","0000000101000","0000000100101","0000000100001","0000000011110","0000000011011","0000000011000","0000000010101","0000000010010","0000000001111","0000000001100","0000000001010","0000000000111","0000000000101","0000000000011","0000000000000","1111111111110","1111111111100","1111111111011","1111111111001","1111111110111","1111111110110","1111111110101"),
("1111111011111","1111111011100","1111111011001","1111111010110","1111111010100","1111111010001","1111111001111","1111111001101","1111111001011","1111111001010","1111111001001","1111111001000","1111111001000","1111111001000","1111111001001","1111111001010","1111111001011","1111111001101","1111111001111","1111111010010","1111111010110","1111111011001","1111111011110","1111111100010","1111111100111","1111111101101","1111111110011","1111111111001","1111111111111","0000000000101","0000000001100","0000000010011","0000000011010","0000000100001","0000000101000","0000000101111","0000000110101","0000000111100","0000001000010","0000001001000","0000001001101","0000001010010","0000001010111","0000001011011","0000001011111","0000001100010","0000001100100","0000001100110","0000001101000","0000001101000","0000001101000","0000001101000","0000001100110","0000001100100","0000001100010","0000001011111","0000001011011","0000001010111","0000001010010","0000001001101","0000001001000","0000001000010","0000000111100","0000000110101","0000000101111","0000000101000","0000000100001","0000000011010","0000000010011","0000000001100","0000000000101","1111111111111","1111111111001","1111111110011","1111111101101","1111111100111","1111111100010","1111111011110","1111111011001","1111111010110","1111111010010","1111111001111","1111111001101","1111111001011","1111111001010","1111111001001","1111111001000","1111111001000","1111111001000","1111111001001","1111111001010","1111111001011","1111111001101","1111111001111","1111111010001","1111111010100","1111111010110","1111111011001","1111111011100","1111111011111"),
("0000000001001","0000000001100","0000000010000","0000000010011","0000000010111","0000000011010","0000000011101","0000000100000","0000000100010","0000000100011","0000000100100","0000000100011","0000000100001","0000000011110","0000000011010","0000000010100","0000000001101","0000000000100","1111111111011","1111111110001","1111111100111","1111111011100","1111111010001","1111111000110","1111110111100","1111110110011","1111110101011","1111110100101","1111110100001","1111110011111","1111110011111","1111110100001","1111110100110","1111110101110","1111110110111","1111111000011","1111111010001","1111111100001","1111111110001","0000000000011","0000000010101","0000000100111","0000000111001","0000001001001","0000001011000","0000001100110","0000001110001","0000001111010","0000001111111","0000010000010","0000010000010","0000001111111","0000001111010","0000001110001","0000001100110","0000001011000","0000001001001","0000000111001","0000000100111","0000000010101","0000000000011","1111111110001","1111111100001","1111111010001","1111111000011","1111110110111","1111110101110","1111110100110","1111110100001","1111110011111","1111110011111","1111110100001","1111110100101","1111110101011","1111110110011","1111110111100","1111111000110","1111111010001","1111111011100","1111111100111","1111111110001","1111111111011","0000000000100","0000000001101","0000000010100","0000000011010","0000000011110","0000000100001","0000000100011","0000000100100","0000000100011","0000000100010","0000000100000","0000000011101","0000000011010","0000000010111","0000000010011","0000000010000","0000000001100","0000000001001"),
("0000000001010","0000000000100","1111111111100","1111111110100","1111111101100","1111111100111","1111111100011","1111111100010","1111111100100","1111111101001","1111111110000","1111111110111","1111111111111","0000000000101","0000000001001","0000000001001","0000000000111","0000000000011","1111111111101","1111111110111","1111111110100","1111111110100","1111111111000","0000000000010","0000000010001","0000000100011","0000000110111","0000001001010","0000001011001","0000001100001","0000001011111","0000001010001","0000000111000","0000000010101","1111111101010","1111110111010","1111110001100","1111101100011","1111101000110","1111100110111","1111100111011","1111101010010","1111101111011","1111110110011","1111111110100","0000000111010","0000001111101","0000010110110","0000011100000","0000011110110","0000011110110","0000011100000","0000010110110","0000001111101","0000000111010","1111111110100","1111110110011","1111101111011","1111101010010","1111100111011","1111100110111","1111101000110","1111101100011","1111110001100","1111110111010","1111111101010","0000000010101","0000000111000","0000001010001","0000001011111","0000001100001","0000001011001","0000001001010","0000000110111","0000000100011","0000000010001","0000000000010","1111111111000","1111111110100","1111111110100","1111111110111","1111111111101","0000000000011","0000000000111","0000000001001","0000000001001","0000000000101","1111111111111","1111111110111","1111111110000","1111111101001","1111111100100","1111111100010","1111111100011","1111111100111","1111111101100","1111111110100","1111111111100","0000000000100","0000000001010"),
("0000000000100","0000000000010","1111111111101","1111111111011","1111111111111","0000000001001","0000000010111","0000000011111","0000000011011","0000000001011","1111111110100","1111111100000","1111111011000","1111111100000","1111111110001","0000000000010","0000000001010","0000000000101","1111111111010","1111111110100","1111111111101","0000000010101","0000000110011","0000001000101","0000000111110","0000000011001","1111111100101","1111110110111","1111110100101","1111110110101","1111111011101","0000000000110","0000000011001","0000000001101","1111111110010","1111111100010","1111111111000","0000000111010","0000010010001","0000011001110","0000011000001","0000001010101","1111110100000","1111011100011","1111001101111","1111010000010","1111100101000","0000000101111","0000100110111","0000111011100","0000111011100","0000100110111","0000000101111","1111100101000","1111010000010","1111001101111","1111011100011","1111110100000","0000001010101","0000011000001","0000011001110","0000010010001","0000000111010","1111111111000","1111111100010","1111111110010","0000000001101","0000000011001","0000000000110","1111111011101","1111110110101","1111110100101","1111110110111","1111111100101","0000000011001","0000000111110","0000001000101","0000000110011","0000000010101","1111111111101","1111111110100","1111111111010","0000000000101","0000000001010","0000000000010","1111111110001","1111111100000","1111111011000","1111111100000","1111111110100","0000000001011","0000000011011","0000000011111","0000000010111","0000000001001","1111111111111","1111111111011","1111111111101","0000000000010","0000000000100"),
("1111111111101","0000000000100","1111111111011","0000000000011","0000000011010","0000000010010","1111111101101","1111111100010","1111111111100","0000000000111","1111111111001","0000000000101","0000000100110","0000000011011","1111111100100","1111111010011","1111111111010","0000000001010","1111111110110","0000000000111","0000000111001","0000000101000","1111111010101","1111110111101","1111111110111","0000000001111","1111111110000","0000000001011","0000001011001","0000000111111","1111110111101","1111110010110","1111111110001","0000000011000","1111111100110","0000000010011","0000010011000","0000001101111","1111110000111","1111100111001","1111111100011","0000000110010","1111111001000","0000000101100","0000110000101","0000100111111","1111001100110","1110010100011","1111101000001","0001101011010","0001101011010","1111101000001","1110010100011","1111001100110","0000100111111","0000110000101","0000000101100","1111111001000","0000000110010","1111111100011","1111100111001","1111110000111","0000001101111","0000010011000","0000000010011","1111111100110","0000000011000","1111111110001","1111110010110","1111110111101","0000000111111","0000001011001","0000000001011","1111111110000","0000000001111","1111111110111","1111110111101","1111111010101","0000000101000","0000000111001","0000000000111","1111111110110","0000000001010","1111111111010","1111111010011","1111111100100","0000000011011","0000000100110","0000000000101","1111111111001","0000000000111","1111111111100","1111111100010","1111111101101","0000000010010","0000000011010","0000000000011","1111111111011","0000000000100","1111111111101"),
("1111111101011","0000000000100","1111111111100","0000000011001","1111111100110","0000000000101","1111111111011","0000000011111","1111111100000","0000000000110","1111111111010","0000000100110","1111111011000","0000000000111","1111111111000","0000000101110","1111111010000","0000000001001","1111111110111","0000000111000","1111111000101","0000000001011","1111111110101","0000001000101","1111110110111","0000000001101","1111111110010","0000001010110","1111110100101","0000000010001","1111111101110","0000001101110","1111110001011","0000000010110","1111111101001","0000010010001","1111101100011","0000000011101","1111111100000","0000011001110","1111100011011","0000000101100","1111111001110","0000101010011","1111001101110","0000001010100","1111110010011","0001101111001","1101000110100","0001011111100","0001011111100","1101000110100","0001101111001","1111110010011","0000001010100","1111001101110","0000101010011","1111111001110","0000000101100","1111100011011","0000011001110","1111111100000","0000000011101","1111101100011","0000010010001","1111111101001","0000000010110","1111110001011","0000001101110","1111111101110","0000000010001","1111110100101","0000001010110","1111111110010","0000000001101","1111110110111","0000001000101","1111111110101","0000000001011","1111111000101","0000000111000","1111111110111","0000000001001","1111111010000","0000000101110","1111111111000","0000000000111","1111111011000","0000000100110","1111111111010","0000000000110","1111111100000","0000000011111","1111111111011","0000000000101","1111111100110","0000000011001","1111111111100","0000000000100","1111111101011"));


-- components 

-- The samples come from the main main 
-- The Coefficents will be here or in the package 

-- serialfilter component 
COMPONENT serial_filter IS 
  GENERIC(
        NUM_OF_COEFFS : NATURAL );
    PORT( 
        clk     : IN STD_LOGIC;
        reset   : IN STD_LOGIC;
        CO      : IN coefficient_type;
        CE      : IN STD_LOGIC;
        sample1 : IN sample;
        sample2 : IN sample;
        Q	      : OUT Multi_Result);
END COMPONENT;

-- signals 
--SIGNAL CE_FIR1,OE_FIR1,CE_FIR2,OE_FIR2: STD_LOGIC; Not used ?? /shwan
SIGNAL Q_FIR1, Q_FIR2 :  Multi_Result;
SIGNAL CO_FIR1,CO_FIR2 : coefficient_type;

SIGNAL start_filter : STD_LOGIC;

BEGIN 
-- component instantiation 
FIR1:  serial_filter 
    GENERIC MAP (
        NUM_OF_COEFFS => NUM_OF_COEFFS)
    PORT MAP(
        clk => clk,
        reset => updated,
        CO => CO_FIR1,
        CE => start_filter,
        sample1 => sample1,
        sample2 => sample2,
        Q => Q_FIR1);
    
FIR2:  serial_filter
    GENERIC MAP (
        NUM_OF_COEFFS => NUM_OF_COEFFS)
    PORT MAP(
        clk => clk,
        reset => updated,
        CO => CO_FIR2,
        CE => start_filter,
        sample1 => sample1,
        sample2 => sample2,
        Q => Q_FIR2);

PROCESS(clk, updated)
    VARIABLE count : NATURAL RANGE 0 TO NUM_OF_COEFFS;
    VARIABLE count_filters : NATURAL RANGE 0 TO NUM_OF_BANDS+1;
    TYPE state_type IS (IDLE, READ_SAMPLE, UPDATE_FILTER, UPDATE_OUTPUT);
    VARIABLE state : state_type;
    VARIABLE Q_sig : Multi_Result_array;
BEGIN

IF clk'EVENT AND clk = '1' THEN
    IF updated = '1' THEN
        state := READ_SAMPLE;
        count := 0;
        count_filters := 0;
        start_filter <= '0';
        done <= '0';
    ELSE
            CASE (state) IS
                WHEN IDLE =>
                    done <= '0';
                WHEN READ_SAMPLE =>
                    next_sample <= '1';
                    start_filter <= '0';
                    sample_nr <= STD_LOGIC_VECTOR(TO_UNSIGNED(count, 7));
                    state := UPDATE_FILTER;
                    
                WHEN UPDATE_FILTER =>
                    next_sample <= '0';
                    CO_FIR1 <= CO(count_filters, count);
                    CO_FIR2 <= CO(count_filters+1, count);
                    start_filter <= '1';
                    IF count < NUM_OF_COEFFS-1 THEN
                        count := count + 1;
                        state := READ_SAMPLE;
                    ELSE
                        count := 0;
                        state := UPDATE_OUTPUT;
                    END IF;
                    
                WHEN UPDATE_OUTPUT =>
                    Q_sig(count_filters) := Q_FIR1;
                    Q_sig(count_filters+1) := Q_FIR2;
                    start_filter <= '0';
                    IF count_filters < NUM_OF_BANDS-2 THEN
                        count_filters := count_filters + 2; -- since we calculate 2 filters at the time
                        state := READ_SAMPLE;
                    ELSE
                        done <= '1';
                        count_filters := 0;
						Q <= Q_sig;
                        state := IDLE;
                    END IF;
            END CASE;
        END IF;
END IF; --clk
END PROCESS;

END ARCHITECTURE;
