-- Description:
-- filterblock_main.vhd
-- Author: Shwan Ciyako,Anandhavel Sakthivel
-- It is still in the implementation phase. 
-- This files adds needed components together to make a filterbank, you are welcome to make changes but make shure to update the whole chain of files that will be affected
--DEMO VERSIOM
-- NO CHANGES ARE ALLOWED IF NOT ANAND IS CONTATED EVEN IF IT IS 6 AM !! 
-- The code is woring fine now by using the updated as trigger to start and oe as the ouput , OE is 
-- updated to one for one cycle as the same time as the Q is putted out, remember it might happen that you catch OE and update your input with the old values 
-- and you need to make sure that some thing like WAIT DATA STate here is implmented to sample this output one clock after the OE goes high. 
-- GOOD LUCK
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_signed.ALL;
USE work.EQ_data_type.ALL;
USE work.EQ_functions.ALL;

ENTITY filterblock_main IS
      GENERIC(
            NUM_BITS_OUT : NATURAL := 13;
            NUM_OF_SAMPLES : NATURAL := 200;
                    NUM_OF_COEFFS : NATURAL := 110;
            NUM_OF_BANDS: NATURAL := 8);
    PORT( 
            clk     : IN STD_LOGIC;
            reset   : IN STD_LOGIC;
            CE      : IN STD_LOGIC;
            sample1 : IN sample;
            sample2 : IN sample;
            updated: IN STD_LOGIC;  -- works as STARTED here no need to add more signals
                RE      : OUT STD_LOGIC;
            OE      : OUT STD_LOGIC; 
            Q       : OUT Multi_Result_array);
END filterblock_main;

ARCHITECTURE  filterblock_main_arch OF filterblock_main IS 
-- constants 
CONSTANT CO:taps_type:=(
("000000000000100101101100","000000000000100101111011","000000000000100110010101","000000000000100110111010","000000000000100111101100","000000000000101000101000","000000000000101001110001","000000000000101011000110","000000000000101100100111","000000000000101110010011","000000000000110000001100","000000000000110010010000","000000000000110100100001","000000000000110110111110","000000000000111001100110","000000000000111100011011","000000000000111111011011","000000000001000010100111","000000000001000101111111","000000000001001001100011","000000000001001101010010","000000000001010001001100","000000000001010101010010","000000000001011001100011","000000000001011101111111","000000000001100010100110","000000000001100111010111","000000000001101100010100","000000000001110001011010","000000000001110110101010","000000000001111100000100","000000000010000001101000","000000000010000111010101","000000000010001101001100","000000000010010011001011","000000000010011001010011","000000000010011111100011","000000000010100101111011","000000000010101100011010","000000000010110011000010","000000000010111001110000","000000000011000000100100","000000000011000111100000","000000000011001110100001","000000000011010101101000","000000000011011100110100","000000000011100100000101","000000000011101011011011","000000000011110010110101","000000000011111010010010","000000000100000001110011","000000000100001001010111","000000000100010000111110","000000000100011000100110","000000000100100000010001","000000000100100111111101","000000000100101111101001","000000000100110111010110","000000000100111111000100","000000000101000110110000","000000000101001110011101","000000000101010110000111","000000000101011101110001","000000000101100101011000","000000000101101100111100","000000000101110100011110","000000000101111011111100","000000000110000011010111","000000000110001010101101","000000000110010001111111","000000000110011001001100","000000000110100000010011","000000000110100111010100","000000000110101110001111","000000000110110101000100","000000000110111011110001","000000000111000010010111","000000000111001000110101","000000000111001111001010","000000000111010101011000","000000000111011011011100","000000000111100001010111","000000000111100111001000","000000000111101100101111","000000000111110010001100","000000000111110111011110","000000000111111100100110","000000001000000001100010","000000001000000110010010","000000001000001010110111","000000001000001111001111","000000001000010011011011","000000001000010111011011","000000001000011011001110","000000001000011110110011","000000001000100010001011","000000001000100101010110","000000001000101000010011","000000001000101011000011","000000001000101101100100","000000001000101111110111","000000001000110001111100","000000001000110011110010","000000001000110101011010","000000001000110110110011","000000001000110111111101","000000001000111000111001","000000001000111001100110","000000001000111010000100","000000001000111010010011"),
("111111111111000000111010","111111111111000011000000","111111111111000100110111","111111111111000110100001","111111111111000111111111","111111111111001001010100","111111111111001010100011","111111111111001011101101","111111111111001100110101","111111111111001101111101","111111111111001111000111","111111111111010000010110","111111111111010001101100","111111111111010011001100","111111111111010100110111","111111111111010110110000","111111111111011000111010","111111111111011011010110","111111111111011110001000","111111111111100001010000","111111111111100100110010","111111111111101000101111","111111111111101101001010","111111111111110010000100","111111111111110111100000","111111111111111101011111","000000000000000100000100","000000000000001011001111","000000000000010011000011","000000000000011011100000","000000000000100100101010","000000000000101110100000","000000000000111001000100","000000000001000100011000","000000000001010000011011","000000000001011101010000","000000000001101010110111","000000000001111001010001","000000000010001000011101","000000000010011000011101","000000000010101001010001","000000000010111010111001","000000000011001101010101","000000000011100000100100","000000000011110100101000","000000000100001001011110","000000000100011111001000","000000000100110101100011","000000000101001100110000","000000000101100100101101","000000000101111101011010","000000000110010110110100","000000000110110000111100","000000000111001011101111","000000000111100111001100","000000001000000011010001","000000001000011111111100","000000001000111101001100","000000001001011010111111","000000001001111001010010","000000001010011000000010","000000001010110111001111","000000001011010110110101","000000001011110110110010","000000001100010111000011","000000001100110111100110","000000001101011000010111","000000001101111001010101","000000001110011010011011","000000001110111011100111","000000001111011100110111","000000001111111110000111","000000010000011111010100","000000010001000000011010","000000010001100001010111","000000010010000010001000","000000010010100010101010","000000010011000010111000","000000010011100010110001","000000010100000010010000","000000010100100001010011","000000010100111111110111","000000010101011101111000","000000010101111011010100","000000010110011000000111","000000010110110100001110","000000010111001111100111","000000010111101010001111","000000011000000100000010","000000011000011100111111","000000011000110101000010","000000011001001100001001","000000011001100010010001","000000011001110111011000","000000011010001011011101","000000011010011110011100","000000011010110000010011","000000011011000001000001","000000011011010000100101","000000011011011110111011","000000011011101100000011","000000011011110111111011","000000011100000010100010","000000011100001011110110","000000011100010011111000","000000011100011010100101","000000011100011111111101","000000011100100011111111","000000011100100110101100","000000011100101000000011"),
("000000000000001000000100","000000000000000001000000","111111111111111001110110","111111111111110010100000","111111111111101010111010","111111111111100010111101","111111111111011010100101","111111111111010001101011","111111111111001000001011","111111111110111110000001","111111111110110011001000","111111111110100111011100","111111111110011010111001","111111111110001101011100","111111111101111111000010","111111111101101111101010","111111111101011111010010","111111111101001101110111","111111111100111011011011","111111111100100111111101","111111111100010011011110","111111111011111101111111","111111111011100111100010","111111111011010000001011","111111111010110111111011","111111111010011110111000","111111111010000101000110","111111111001101010101011","111111111001001111101011","111111111000110100001111","111111111000011000011101","111111110111111100011100","111111110111100000010110","111111110111000100010010","111111110110101000011010","111111110110001100110111","111111110101110001110100","111111110101010111011010","111111110100111101110100","111111110100100101001101","111111110100001101101111","111111110011110111100110","111111110011100010111101","111111110011001111111110","111111110010111110110101","111111110010101111101100","111111110010100010101101","111111110010011000000100","111111110010001111111001","111111110010001010010111","111111110010000111100110","111111110010000111101111","111111110010001010111010","111111110010010001001111","111111110010011010110011","111111110010100111101110","111111110010111000000100","111111110011001011111001","111111110011100011010010","111111110011111110010000","111111110100011100110110","111111110100111111000011","111111110101100100111001","111111110110001110010110","111111110110111011010111","111111110111101011111001","111111111000011111111000","111111111001010111001111","111111111010010001111000","111111111011001111101011","111111111100010000011111","111111111101010100001101","111111111110011010101001","111111111111100011101000","000000000000101110111111","000000000001111100100001","000000000011001100000000","000000000100011101001110","000000000101101111111101","000000000111000011111011","000000001000011000111010","000000001001101110101001","000000001011000100110111","000000001100011011010010","000000001101110001101000","000000001111000111101000","000000010000011100111111","000000010001110001011100","000000010011000100101100","000000010100010110011101","000000010101100110011110","000000010110110100011100","000000011000000000000111","000000011001001001001101","000000011010001111011110","000000011011010010101011","000000011100010010100011","000000011101001110111001","000000011110000111011110","000000011110111100000110","000000011111101100100011","000000100000011000101100","000000100001000000010110","000000100001100011010111","000000100010000001100111","000000100010011011000000","000000100010101111011011","000000100010111110110100","000000100011001001000110","000000100011001110010000"),
("000000000000100010011001","000000000000101011000101","000000000000110011111101","000000000000111101001000","000000000001000110101001","000000000001010000100100","000000000001011010111100","000000000001100101110011","000000000001110001001100","000000000001111101000111","000000000010001001100011","000000000010010110011111","000000000010100011111000","000000000010110001101010","000000000010111111110001","000000000011001110000101","000000000011011100011111","000000000011101010110110","000000000011111001000000","000000000100000110110001","000000000100010011111101","000000000100100000010111","000000000100101011101111","000000000100110101111000","000000000100111110100010","000000000101000101011100","000000000101001010010111","000000000101001101000011","000000000101001101001111","000000000101001010101011","000000000101000101001001","000000000100111100011010","000000000100110000010001","000000000100100000100011","000000000100001101000011","000000000011110101101010","000000000011011010010000","000000000010111010110000","000000000010010111001000","000000000001101111010110","000000000001000011011100","000000000000010011100000","111111111111011111101000","111111111110100111111101","111111111101101100101110","111111111100101110001000","111111111011101100011110","111111111010101000000101","111111111001100001010101","111111111000011000101000","111111110111001110011001","111111110110000011001000","111111110100110111010101","111111110011101011100011","111111110010100000010110","111111110001010110010011","111111110000001110000010","111111101111001000001000","111111101110000101001101","111111101101000101111011","111111101100001010110110","111111101011010100101000","111111101010100011110101","111111101001111001000001","111111101001010100110001","111111101000110111100100","111111101000100001111001","111111101000010100001100","111111101000001110110110","111111101000010010001100","111111101000011110011111","111111101000110011111111","111111101001010010110110","111111101001111011001000","111111101010101100111001","111111101011101000000101","111111101100101100100100","111111101101111010001011","111111101111010000101001","111111110000101111101010","111111110010010110110011","111111110100000101101000","111111110101111011100101","111111110111111000000101","111111111001111010011111","111111111100000010000100","111111111110001110000101","000000000000011101101110","000000000010110000001001","000000000101000100011111","000000000111011001110101","000000001001101111010010","000000001100000011111000","000000001110010110101101","000000010000100110110011","000000010010110011001111","000000010100111011000111","000000010110111101100010","000000011000111001101000","000000011010101110100100","000000011100011011100101","000000011101111111111011","000000011111011010111010","000000100000101011111100","000000100001110010011101","000000100010101101111111","000000100011011110000110","000000100100000010011110","000000100100011010110111","000000100100100111000110"),
("111111111111011011011101","111111111111011011000010","111111111111011011001001","111111111111011011110001","111111111111011100111000","111111111111011110011100","111111111111100000011101","111111111111100010111000","111111111111100101101011","111111111111101000110001","111111111111101100000111","111111111111101111100110","111111111111110011001000","111111111111110110100011","111111111111111001101111","111111111111111100100001","111111111111111110101101","000000000000000000000111","000000000000000000100100","111111111111111111110110","111111111111111101110101","111111111111111010010101","111111111111110101010001","111111111111101110100011","111111111111100110001011","111111111111011100001100","111111111111010000101110","111111111111000011111101","111111111110110110001011","111111111110100111110001","111111111110011001001001","111111111110001010110111","111111111101111101100001","111111111101110001110001","111111111101101000010100","111111111101100001111011","111111111101011111010110","111111111101100001010101","111111111101101000100110","111111111101110101110100","111111111110001001100010","111111111110100100001111","111111111111000110001111","111111111111101111101101","000000000000100000101001","000000000001011000110011","000000000010010111110001","000000000011011100110111","000000000100100111001101","000000000101110101101010","000000000111000110111000","000000001000011001010101","000000001001101011010001","000000001010111010110010","000000001100000101110111","000000001101001010011000","000000001110000110001110","000000001110110111001101","000000001111011011010001","000000001111110000011101","000000001111110100111100","000000001111100111001010","000000001111000101110100","000000001110001111111011","000000001101000100111001","000000001011100100100000","000000001001101110111111","000000000111100101000100","000000000101000111111001","000000000010011001000110","111111111111011010110010","111111111100001111100000","111111111000111010001101","111111110101011110001111","111111110001111111001111","111111101110100001000111","111111101011000111111101","111111100111110111111101","111111100100110101010110","111111100010000100010010","111111011111101000110011","111111011101100110101000","111111011100000001010000","111111011010111011101011","111111011010011000011110","111111011010011001100111","111111011011000000011110","111111011100001101110011","111111011110000001100101","111111100000011011001001","111111100011011001000010","111111100110111001001001","111111101010111000101000","111111101111010100000001","111111110100000111001111","111111111001001101101100","111111111110100010010011","000000000011111111101010","000000001001100000000110","000000001110111101110011","000000010100010010111000","000000011001011001100011","000000011110001100001101","000000100010100101100001","000000100110100000100110","000000101001111001000000","000000101100101010111100","000000101110110011001111","000000110000001111011111","000000110000111110000001"),
("000000000000110011111100","000000000000110110001011","000000000000110101010110","000000000000110001001100","000000000000101001101100","000000000000011110111110","000000000000010001011011","000000000000000001101011","111111111111110000100000","111111111111011110111100","111111111111001110000101","111111111110111111001000","111111111110110011001101","111111111110101011010100","111111111110101000001110","111111111110101010010110","111111111110110001101001","111111111110111101101010","111111111111001101011011","111111111111011111100110","111111111111110010011101","000000000000000100001010","000000000000010010110110","000000000000011100111010","000000000000100001001011","000000000000011111000011","000000000000010110110010","000000000000001001011010","111111111111111000110001","111111111111100111011110","111111111111011000100110","111111111111001111011001","111111111111001111000001","111111111111011010000101","111111111111110010010000","000000000000011000000010","000000000001001010011001","000000000010000110110010","000000000011001001000111","000000000100001100000000","000000000101001001001010","000000000101111001111001","000000000110010111101101","000000000110011101000000","000000000110000101101100","000000000101001111110001","000000000011111011101101","000000000010001100101011","000000000000001000011100","111111111101110111001001","111111111011100010101000","111111111001010101110010","111111110111011011100000","111111110101111101101110","111111110101000100011101","111111110100110100110110","111111110101010000100110","111111110110010101100110","111111110111111101111001","111111111010000000001000","111111111100010000001111","111111111110100000100110","000000000000100011010010","000000000010001011100100","000000000011001111001111","000000000011100111111011","000000000011010100000010","000000000010010111010000","000000000000111010100110","111111111111001011110111","111111111101011100100001","111111111100000000010000","111111111011001010111101","111111111011001110101011","111111111100011001011100","111111111110110011010110","000000000010011101000011","000000000111001110101111","000000001100110111111101","000000010011000000000110","000000011001000111110110","000000011110101011010001","000000100011000100100100","000000100101101111001100","000000100110001011010001","000000100100000000110011","000000011111000010011010","000000010111001111101000","000000001100110101111110","000000000000010001010000","111111110010001010100000","111111100011010101110111","111111010100101111011010","111111000111010111001010","111110111100001100011111","111110110100001001010111","111110101111111101110000","111110110000001011011110","111110110101000011000100","111110111110100001101100","111111001100010000100010","111111011101100101100000","111111110001100101100110","000000000111001000011010","000000011100111100110100","000000110001101110010101","000001000100001010111111","000001010011001000111001","000001011101101011100010","000001100011000111111111"),
("111111111111001010011100","111111111111010001001001","111111111111100001000100","111111111111110100010011","000000000000000100010100","000000000000001100001010","000000000000001010010001","000000000000000001000111","111111111111110110011110","111111111111110001011100","111111111111110111101010","000000000000001010111000","000000000000100111100000","000000000001000101000100","000000000001011000101101","000000000001011000101101","000000000001000000011100","000000000000010010110000","111111111111011010000010","111111111110100101100010","111111111110000100011001","111111111110000000011010","111111111110011010000100","111111111111000111101111","111111111111111000110011","000000000000011011100001","000000000000100100001101","000000000000010010010011","111111111111110001101111","111111111111010111000101","111111111111010111101011","000000000000000000011010","000000000001001110100111","000000000010101110010001","000000000011111111000001","000000000100011110110011","000000000011110110100110","000000000010000100110001","111111111111100000011011","111111111100110100000110","111111111010110000011110","111111111001111011101010","111111111010100011001011","111111111100010101110100","111111111110101000110100","000000000000100111000110","000000000001100101010110","000000000001010011101011","000000000000000101101000","111111111110101100011111","111111111110000100111010","111111111110111110001000","000000000001100011101001","000000000101010010110110","000000001001000001110000","000000001011010110000100","000000001011000101011110","000000000111110011100001","000000000010000001101111","111111111011001010001111","111111110101000101001100","111111110001100001001011","111111110001011100001011","111111110100101011110101","111111111001111111000110","111111111111011010000001","000000000011000011011000","000000000011110011011111","000000000001110010100010","111111111110011001011010","111111111011110010010100","111111111100000010110101","000000000000010010010101","000000001000000011000101","000000010001001110110001","000000011000101011101001","000000011011001111111111","000000010110111101100010","000000001011111001011000","111111111100011001011100","111111101100011110101101","111111100000100101100110","111111011100000110000010","111111100000000101000110","111111101010110110100000","111111111000011100101101","000000000100000000101111","000000001001100101011100","000000000111101101010101","000000000000001011100001","111111110111101000000000","111111110011111010001001","111111111001110111000001","000000001011000101010001","000000100100101010110110","000000111111011010010001","000001010001100110111101","000001010010000100110100","000000111011011010010001","000000001110011111101000","111111010011010000011111","111110010111010011000011","111101101010100010111110","111101011010110111001100","111101101111110011110111","111110100111111011101000","111111111000011011001110","000001001111011110101011","000010011000101100011100","000011000010011010000100"),
("000000000000110000011011","000000000000101110001010","111111111111111110110110","111111111111001110111011","111111111111001100110100","111111111111110001101000","000000000000001100010001","000000000000000010001110","111111111111110010000100","000000000000000111101101","000000000000111001010000","000000000001001000111011","000000000000010010010110","111111111111000010011001","111111111110101001001111","111111111111011001000100","000000000000001111000011","000000000000001011111011","111111111111101010111100","111111111111111101001011","000000000001010000001011","000000000010000101001010","000000000001000001010101","111111111110110000000000","111111111101100001011110","111111111110011110010100","000000000000001010111100","000000000000100000100001","111111111111100101001010","111111111111100101110001","000000000001100111111001","000000000011100110011000","000000000010100100011110","111111111110101111110010","111111111011110100111101","111111111100101010101110","111111111111101100111110","000000000001000001110100","111111111111101011001111","111111111110111101110101","000000000001101110001011","000000000101100101100001","000000000101010010010100","111111111111100101001011","111111111001110000010001","111111111001100111111111","111111111110010110100010","000000000001101000110001","000000000000001011010000","111111111110001001111111","000000000001001111111011","000000000111110001001010","000000001001011100001011","000000000001111101100100","111111110111101111110011","111111110101000011001011","111111111011011100000001","000000000010000000011010","000000000001010011011010","111111111101011000011010","111111111111111100110111","000000001001101111111000","000000001111001111001010","000000000110110010001010","111111110110100001111110","111111101110101011110001","111111110101111111000110","000000000001011111001111","000000000011001110111001","111111111101000001001111","111111111101101000110110","000000001011000011110110","000000010110111110011100","000000001111010111000100","111111110111001110010111","111111100110001000000101","111111101100010111001011","111111111110110110111000","000000000110000101011111","111111111101101001010010","111111111010000110000011","000000001011001100000111","000000100001100111110110","000000011110011011001010","111111111011110111000110","111111011010000110011100","111111011010101111000110","111111110111010100110000","000000001010000101001111","000000000000010111000001","111111110100100110001100","000000001001010111100110","000000110011001111000000","000000111101000010010101","000000001010010011011011","111111000100101111001010","111110110010010111011101","111111100000011111001010","000000010000101000110011","000000001001011001101111","111111101000011011111100","000000000010010110111101","000001101000001100010101","000010101101000100101001","000001010000000111110011","111101100111000101100011","111010111010101111010000","111100001111001010111001","000001001000110111100111","000101100100100010110100")
);


-- components 

-- The samples come from the main main 
-- The Coefficents will be here or in the package 

-- serialfilter component 
COMPONENT serial_filter IS 
  GENERIC(
        NUM_BITS_OUT : NATURAL := 37;
        NUM_OF_COEFFS : NATURAL := 110);
PORT( 
        clk     : IN STD_LOGIC;
        reset   : IN STD_LOGIC;
        CO      : IN coefficient_type;
        CE      : IN STD_LOGIC;
        sample1 : IN sample;
        sample2 : IN sample;
        updated : IN STD_LOGIC;
        OE      : OUT STD_LOGIC;
        Q        : OUT Multi_Result);
    --  Q       : OUT STD_LOGIC_VECTOR(NUM_BITS_OUT-1 DOWNTO 0));
END COMPONENT;


-- signals 
SIGNAL OE_FIR1,OE_FIR2: STD_LOGIC; --CE_FIR1,CE_FIR2,
SIGNAL Q_FIR1,Q_FIR2 :  Multi_Result;
SIGNAL CO_FIR1,CO_FIR2 : coefficient_type;

TYPE state_type_Filter_Bank IS ( WAIT_SAMPLE, COMPUTE_DATA, WAIT_DATA, OUTPUT_DATA);
SIGNAL STATE : state_type_Filter_Bank;
SIGNAL Q_sig: Multi_Result_array;
SIGNAL startfilters: STD_LOGIC;
BEGIN 
-- component instantiation 
FIR1: serial_filter PORT MAP(clk,reset,CO_FIR1,CE,sample1,sample2,startfilters,OE_FIR1,Q_FIR1);
FIR2:  serial_filter PORT MAP(clk,reset,CO_FIR2,CE,sample1,sample2,startfilters,OE_FIR2,Q_FIR2);

---------- Process updating the current state -----------
--update_state: PROCESS ( clk )
--BEGIN
--    IF clk'EVENT and clk = '1' THEN
--        state <= next_state;
--    END IF;
--END PROCESS update_state;

PROCESS(clk,reset,CE,sample1,sample2,updated)
----------Variables -------------------------------------

    VARIABLE count : NATURAL RANGE 0 TO NUM_OF_COEFFS;
    VARIABLE count_filters : NATURAL RANGE 0 TO NUM_OF_BANDS;
    
---------------------------------------------------------
BEGIN

IF clk'EVENT AND clk = '1' THEN
        -- Synchronous reset
        IF reset ='1' THEN 
                FOR k IN 1 TO 8 LOOP
                Q(k) <= (OTHERS => '0');
                          Q_sig(k) <= (OTHERS => '0');
                END LOOP;
                          count := 0;
                          count_filters:=1;
                OE    <= '0';
                STATE <= WAIT_SAMPLE ;
                 RE<= '0';

        ELSIF CE = '1' THEN -- slow clock
        
        CASE STATE IS 
        
          WHEN WAIT_SAMPLE => 
                OE <= '0';
                
                  IF UPDATED = '1' THEN
                     RE <= '1'; 
                     startfilters <='1';
                     STATE <= COMPUTE_DATA ; 
                END IF ; --updated
            
          WHEN COMPUTE_DATA =>
            -- same CE for the filters and the buffer will result in one value per CE moved from buffers to the filters 
           
                 IF count_filters < ((NUM_OF_BANDS/2)+1) then -- 4 filters right now are serially implemented can be changed
            
                    IF count < NUM_OF_COEFFS then 
                     OE<='0';
                     -- move this ?
                 startfilters <='0';
                       CO_FIR1 <= CO(count_filters,count+1);
                       CO_FIR2 <= CO(count_filters+((NUM_OF_BANDS/2)),count+1); -- this start from 4 right/anand
                       count := count +1;
                       ELSE 
                       count := 0;
                       state <= WAIT_DATA;
                   -- this is a test 
                       --Q_sig(count_filters) <= Q_FIR1;
                       --Q_sig(count_filters+(NUM_OF_BANDS/2)) <= Q_FIR2;
                       
                       END IF; -- count
                     ELSE 
                       state <= OUTPUT_DATA;
            END IF; 
  
            WHEN WAIT_DATA => 
			IF OE_FIR1 = '1' then
					Q_sig(count_filters) <= Q_FIR1;
                    Q_sig(count_filters+(NUM_OF_BANDS/2)) <= Q_FIR2;
					IF count_filters < ((NUM_OF_BANDS/2)) then		
					startfilters <='1';
                    STATE <= COMPUTE_DATA;
					count_filters := count_filters + 1 ;
					ELSE 
					STATE <= OUTPUT_DATA;
					END IF;
					
			ELSE 
			state <= WAIT_DATA;
			END IF;
            WHEN OUTPUT_DATA =>
             --  convert to state ELSE -- update the output after 4 cycles ie the 8 filters are done
                   Q<= Q_sig;  
                     OE <='1';
                     count := 0;
                     count_filters := 1;
                     startfilters <='0';
                     STATE <= WAIT_SAMPLE;
                     RE<= '0';
                
                
            END CASE;
        
        
        END IF; --reset 
END IF; --clk
End process;

END ARCHITECTURE;
